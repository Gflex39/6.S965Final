module inverse_quantizer(
    input wire clk_in,
    input wire rst_in,
    input wire [95:0] column_in,
    input wire valid_in,

    output logic [95:0] column_out,
    output logic valid_out
);
    logic [2:0] counter;

    logic signed [11:0] c [7:0];
    logic signed [11:0] o [7:0];

    assign c[0] = column_in[11: 0];
    assign c[1] = column_in[23:12];
    assign c[2] = column_in[35:24];
    assign c[3] = column_in[47:36];
    assign c[4] = column_in[59:48];
    assign c[5] = column_in[71:60];
    assign c[6] = column_in[83:72];
    assign c[7] = column_in[95:84];

    assign column_out[11: 0] = o[0];
    assign column_out[23:12] = o[1];
    assign column_out[35:24] = o[2];
    assign column_out[47:36] = o[3];
    assign column_out[59:48] = o[4];
    assign column_out[71:60] = o[5];
    assign column_out[83:72] = o[6];
    assign column_out[95:84] = o[7];

    always_ff @(posedge clk_in) begin
        if (rst_in) begin
            counter <= 0;
            valid_out <= 0;
            for (integer i = 0; i < 8; i = i + 1) begin
                o[i] <= 0;
            end
        end else if (valid_in) begin
            counter <= counter + 1;
            valid_out <= 1;
            case (counter)
                3'd0: begin
                    /* 016 */ o[0] <= (c[0]<<<4);
                    /* 012 */ o[1] <= (c[1]<<<3)+(c[1]<<<2);
                    /* 014 */ o[2] <= (c[2]<<<3)+(c[2]<<<2)+(c[2]<<<1);
                    /* 014 */ o[3] <= (c[3]<<<3)+(c[3]<<<2)+(c[3]<<<1);
                    /* 018 */ o[4] <= (c[4]<<<4)+(c[4]<<<1);
                    /* 024 */ o[5] <= (c[5]<<<4)+(c[5]<<<3);
                    /* 049 */ o[6] <= (c[6]<<<5)+(c[6]<<<4)+c[6];
                    /* 072 */ o[7] <= (c[7]<<<6)+(c[7]<<<3);
                end
                3'd1: begin
                    /* 011 */ o[0] <= (c[0]<<<3)+(c[0]<<<1)+c[0];
                    /* 012 */ o[1] <= (c[1]<<<3)+(c[1]<<<2);
                    /* 013 */ o[2] <= (c[2]<<<3)+(c[2]<<<2)+c[2];
                    /* 017 */ o[3] <= (c[3]<<<4)+c[3];
                    /* 022 */ o[4] <= (c[4]<<<4)+(c[4]<<<2)+(c[4]<<<1);
                    /* 035 */ o[5] <= (c[5]<<<5)+(c[5]<<<1)+c[5];
                    /* 064 */ o[6] <= (c[6]<<<6);
                    /* 092 */ o[7] <= (c[7]<<<6)+(c[7]<<<4)+(c[7]<<<3)+(c[7]<<<2);
                end
                3'd2: begin
                    /* 010 */ o[0] <= (c[0]<<<3)+(c[0]<<<1);
                    /* 014 */ o[1] <= (c[1]<<<3)+(c[1]<<<2)+(c[1]<<<1);
                    /* 016 */ o[2] <= (c[2]<<<4);
                    /* 022 */ o[3] <= (c[3]<<<4)+(c[3]<<<2)+(c[3]<<<1);
                    /* 037 */ o[4] <= (c[4]<<<5)+(c[4]<<<2)+c[4];
                    /* 055 */ o[5] <= (c[5]<<<5)+(c[5]<<<4)+(c[5]<<<2)+(c[5]<<<1)+c[5];
                    /* 078 */ o[6] <= (c[6]<<<6)+(c[6]<<<3)+(c[6]<<<2)+(c[6]<<<1);
                    /* 095 */ o[7] <= (c[7]<<<6)+(c[7]<<<4)+(c[7]<<<3)+(c[7]<<<2)+(c[7]<<<1)+c[7];
                end
                3'd3: begin
                    /* 016 */ o[0] <= (c[0]<<<4);
                    /* 019 */ o[1] <= (c[1]<<<4)+(c[1]<<<1)+c[1];
                    /* 024 */ o[2] <= (c[2]<<<4)+(c[2]<<<3);
                    /* 029 */ o[3] <= (c[3]<<<4)+(c[3]<<<3)+(c[3]<<<2)+c[3];
                    /* 056 */ o[4] <= (c[4]<<<5)+(c[4]<<<4)+(c[4]<<<3);
                    /* 064 */ o[5] <= (c[5]<<<6);
                    /* 087 */ o[6] <= (c[6]<<<6)+(c[6]<<<4)+(c[6]<<<2)+(c[6]<<<1)+c[6];
                    /* 098 */ o[7] <= (c[7]<<<6)+(c[7]<<<5)+(c[7]<<<1);
                end
                3'd4: begin
                    /* 024 */ o[0] <= (c[0]<<<4)+(c[0]<<<3);
                    /* 026 */ o[1] <= (c[1]<<<4)+(c[1]<<<3)+(c[1]<<<1);
                    /* 040 */ o[2] <= (c[2]<<<5)+(c[2]<<<3);
                    /* 051 */ o[3] <= (c[3]<<<5)+(c[3]<<<4)+(c[3]<<<1)+c[3];
                    /* 068 */ o[4] <= (c[4]<<<6)+(c[4]<<<2);
                    /* 081 */ o[5] <= (c[5]<<<6)+(c[5]<<<4)+c[5];
                    /* 103 */ o[6] <= (c[6]<<<6)+(c[6]<<<5)+(c[6]<<<2)+(c[6]<<<1)+c[6];
                    /* 112 */ o[7] <= (c[7]<<<6)+(c[7]<<<5)+(c[7]<<<4);
                end
                3'd5: begin
                    /* 040 */ o[0] <= (c[0]<<<5)+(c[0]<<<3);
                    /* 058 */ o[1] <= (c[1]<<<5)+(c[1]<<<4)+(c[1]<<<3)+(c[1]<<<1);
                    /* 057 */ o[2] <= (c[2]<<<5)+(c[2]<<<4)+(c[2]<<<3)+c[2];
                    /* 087 */ o[3] <= (c[3]<<<6)+(c[3]<<<4)+(c[3]<<<2)+(c[3]<<<1)+c[3]; // 64+16+4+2+1
                    /* 109 */ o[4] <= (c[4]<<<6)+(c[4]<<<5)+(c[4]<<<3)+(c[4]<<<2)+c[4]; // 64+32+8+4+1
                    /* 104 */ o[5] <= (c[5]<<<6)+(c[5]<<<5)+(c[5]<<<3); // 64+32+8
                    /* 121 */ o[6] <= (c[6]<<<6)+(c[6]<<<5)+(c[6]<<<4)+(c[6]<<<3)+c[6]; // 64+32+16+8+1
                    /* 100 */ o[7] <= (c[7]<<<6)+(c[7]<<<5)+(c[7]<<<2); // 64+32+4
                end
                3'd6: begin
                    /* 051 */ o[0] <= (c[0]<<<5)+(c[0]<<<4)+(c[0]<<<1)+c[0]; // 32+16+2+1 = 51
                    /* 060 */ o[1] <= (c[1]<<<5)+(c[1]<<<4)+(c[1]<<<3)+(c[1]<<<2); // 32+16+8+4 = 60
                    /* 069 */ o[2] <= (c[2]<<<6)+(c[2]<<<2)+c[2]; // 64+4+1 = 69
                    /* 080 */ o[3] <= (c[3]<<<6)+(c[3]<<<4); // 64+16 = 80
                    /* 103 */ o[4] <= (c[4]<<<6)+(c[4]<<<5)+(c[4]<<<2)+(c[4]<<<1)+c[4]; // 64+32+4+2+1 = 103
                    /* 113 */ o[5] <= (c[5]<<<6)+(c[5]<<<5)+(c[5]<<<4)+c[5]; // 64+32+16+1 = 113
                    /* 120 */ o[6] <= (c[6]<<<6)+(c[6]<<<5)+(c[6]<<<4)+(c[6]<<<3); // 64+32+16+8 = 120
                    /* 103 */ o[7] <= (c[7]<<<6)+(c[7]<<<5)+(c[7]<<<2)+(c[7]<<<1)+c[7];  // 64+32+4+2+1 = 103
                end
                3'd7: begin
                    /* 061 */ o[0] <= (c[0]<<<5)+(c[0]<<<4)+(c[0]<<<3)+(c[0]<<<2)+c[0]; // 32+16+8+4+1 = 61
                    /* 055 */ o[1] <= (c[1]<<<5)+(c[1]<<<4)+(c[1]<<<2)+(c[1]<<<1)+c[1]; // 32+16+4+2+1 = 55
                    /* 056 */ o[2] <= (c[2]<<<5)+(c[2]<<<4)+(c[2]<<<3); // 32+16+8 = 56
                    /* 062 */ o[3] <= (c[3]<<<5)+(c[3]<<<4)+(c[3]<<<3)+(c[3]<<<2)+(c[3]<<<1); // 32+16+8+4+2 = 62
                    /* 077 */ o[4] <= (c[4]<<<6)+(c[4]<<<3)+(c[4]<<<2)+c[4]; // 64+8+4+1 = 77
                    /* 092 */ o[5] <= (c[5]<<<6)+(c[5]<<<4)+(c[5]<<<3)+(c[5]<<2); // 64+16+8+4 = 92
                    /* 101 */ o[6] <= (c[6]<<<6)+(c[6]<<<5)+(c[6]<<<2)+c[6]; // 64+32+4+1 = 101
                    /* 099 */ o[7] <= (c[7]<<<6)+(c[7]<<<5)+(c[7]<<<1)+c[7]; // 64+32+2+1 = 99
                end
            endcase
        end else begin
            valid_out <= 0;
            o[0] <= 0;
            o[1] <= 0;
            o[2] <= 0;
            o[3] <= 0;
            o[4] <= 0;
            o[5] <= 0;
            o[6] <= 0;
            o[7] <= 0;
        end
    end

endmodule