`timescale 1ns / 1ps
`default_nettype none

module zigzag_decoder(
    input wire clk_in,
    input wire rst_in,
    input wire signed [11:0] value_in,
    input wire [4:0] run_in,
    input wire dc_in,
    input wire valid_in
);
endmodule